`timescale 1ns / 1ps

module Data_mem(
    input           CLK,    // ���� �������������
    input   [31:0]   A,     // 32-������ �������� ����
    input   [31:0]  WD,    // 32-������ ���� ������ ��� ������
    input           WE,     // ������ ���������� �� ������
    output [31:0]  RD      // 31-������ ����� ��������� ������
);

  reg [31:0] RAM [0:255];  // ������� ������ � 256-� 32-������� ��������
  
  initial $readmemb("mem.mem", RAM);

  // ������
   assign RD = RAM[A[9:2]];     // ���������� � ������ RD ������ ������ �� ������ A[9:2]

  // ������
  always @ (posedge CLK)  // ������ ���, ����� ���������� ����� CLK
    if (WE)               // ���� ������ WE == 1
      RAM[A[9:2]] <= WD;  // � ������ �� ������ A[9:2] ����� �������� ������ WD

endmodule
